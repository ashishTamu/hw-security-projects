module StraightPBox()
endmodule
