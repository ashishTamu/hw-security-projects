module InitialPermutation()
endmodule
