module Encryption()
endmodule
