library ieee;
use ieee.std_logic_1164.all;
entity scan_chain is port
(
scan_clk : in std_logic;
reset : in std_logic;
test_enable : in std_logic;
ShiftDR : in std_logic;
UpdateDR : in std_logic;
CaptureDR : in std_logic;
scan_in : in std_logic;
li_in,ri_in : in std_logic_vector(1 to 32);
lo_in,ro_in : in std_logic_vector(1 to 32);
li_dataout,ri_dataout: out std_logic_vector(1 to 32);
lo_dataout,ro_dataout : out std_logic_vector(1 to 32);
scan_out : out std_logic
);
end scan_chain;
architecture behaviour of scan_chain is
signal li_1,li_2,li_3,li_4,li_5,li_6,li_7,li_8,li_9,li_10,li_11,li_12,li_13,li_14,li_15,li_16,li_17,li_18,li_19,li_20,li_21,li_22,li_23,li_24,li_25,li_26,li_27,li_28,li_29,li_30,li_31,li_32: std_logic;--_vector (1 to 1);
signal ri_1,ri_2,ri_3,ri_4,ri_5,ri_6,ri_7,ri_8,ri_9,ri_10,ri_11,ri_12,ri_13,ri_14,ri_15,ri_16,ri_17,ri_18,ri_19,ri_20,ri_21,ri_22,ri_23,ri_24,ri_25,ri_26,ri_27,ri_28,ri_29,ri_30,ri_31,ri_32: std_logic;--_vector (1 to 1);
signal lo_1,lo_2,lo_3,lo_4,lo_5,lo_6,lo_7,lo_8,lo_9,lo_10,lo_11,lo_12,lo_13,lo_14,lo_15,lo_16,lo_17,lo_18,lo_19,lo_20,lo_21,lo_22,lo_23,lo_24,lo_25,lo_26,lo_27,lo_28,lo_29,lo_30,lo_31,lo_32: std_logic;--_vector (1 to 1);
signal ro_1,ro_2,ro_3,ro_4,ro_5,ro_6,ro_7,ro_8,ro_9,ro_10,ro_11,ro_12,ro_13,ro_14,ro_15,ro_16,ro_17,ro_18,ro_19,ro_20,ro_21,ro_22,ro_23,ro_24,ro_25,ro_26,ro_27,ro_28,ro_29,ro_30,ro_31,ro_32: std_logic;--_vector (1 to 1);
signal li_scanout_1,li_scanout_2,li_scanout_3,li_scanout_4,li_scanout_5,li_scanout_6,li_scanout_7,li_scanout_8,li_scanout_9,li_scanout_10,li_scanout_11,li_scanout_12,li_scanout_13,li_scanout_14,li_scanout_15,li_scanout_16,li_scanout_17,li_scanout_18,li_scanout_19,li_scanout_20,li_scanout_21,li_scanout_22,li_scanout_23,li_scanout_24,li_scanout_25,li_scanout_26,li_scanout_27,li_scanout_28,li_scanout_29,li_scanout_30,li_scanout_31,li_scanout_32: std_logic;--_vector (1 to 1);
signal ri_scanout_1,ri_scanout_2,ri_scanout_3,ri_scanout_4,ri_scanout_5,ri_scanout_6,ri_scanout_7,ri_scanout_8,ri_scanout_9,ri_scanout_10,ri_scanout_11,ri_scanout_12,ri_scanout_13,ri_scanout_14,ri_scanout_15,ri_scanout_16,ri_scanout_17,ri_scanout_18,ri_scanout_19,ri_scanout_20,ri_scanout_21,ri_scanout_22,ri_scanout_23,ri_scanout_24,ri_scanout_25,ri_scanout_26,ri_scanout_27,ri_scanout_28,ri_scanout_29,ri_scanout_30,ri_scanout_31,ri_scanout_32: std_logic;--_vector (1 to 1);
signal lo_scanout_1,lo_scanout_2,lo_scanout_3,lo_scanout_4,lo_scanout_5,lo_scanout_6,lo_scanout_7,lo_scanout_8,lo_scanout_9,lo_scanout_10,lo_scanout_11,lo_scanout_12,lo_scanout_13,lo_scanout_14,lo_scanout_15,lo_scanout_16,lo_scanout_17,lo_scanout_18,lo_scanout_19,lo_scanout_20,lo_scanout_21,lo_scanout_22,lo_scanout_23,lo_scanout_24,lo_scanout_25,lo_scanout_26,lo_scanout_27,lo_scanout_28,lo_scanout_29,lo_scanout_30,lo_scanout_31,lo_scanout_32: std_logic;--_vector (1 to 1);
signal ro_scanout_1,ro_scanout_2,ro_scanout_3,ro_scanout_4,ro_scanout_5,ro_scanout_6,ro_scanout_7,ro_scanout_8,ro_scanout_9,ro_scanout_10,ro_scanout_11,ro_scanout_12,ro_scanout_13,ro_scanout_14,ro_scanout_15,ro_scanout_16,ro_scanout_17,ro_scanout_18,ro_scanout_19,ro_scanout_20,ro_scanout_21,ro_scanout_22,ro_scanout_23,ro_scanout_24,ro_scanout_25,ro_scanout_26,ro_scanout_27,ro_scanout_28,ro_scanout_29,ro_scanout_30,ro_scanout_31,ro_scanout_32: std_logic;--_vector (1 to 1);
signal li_dataout_1,li_dataout_2,li_dataout_3,li_dataout_4,li_dataout_5,li_dataout_6,li_dataout_7,li_dataout_8,li_dataout_9,li_dataout_10,li_dataout_11,li_dataout_12,li_dataout_13,li_dataout_14,li_dataout_15,li_dataout_16,li_dataout_17,li_dataout_18,li_dataout_19,li_dataout_20,li_dataout_21,li_dataout_22,li_dataout_23,li_dataout_24,li_dataout_25,li_dataout_26,li_dataout_27,li_dataout_28,li_dataout_29,li_dataout_30,li_dataout_31,li_dataout_32: std_logic;--_vector (1 to 1);
signal ri_dataout_1,ri_dataout_2,ri_dataout_3,ri_dataout_4,ri_dataout_5,ri_dataout_6,ri_dataout_7,ri_dataout_8,ri_dataout_9,ri_dataout_10,ri_dataout_11,ri_dataout_12,ri_dataout_13,ri_dataout_14,ri_dataout_15,ri_dataout_16,ri_dataout_17,ri_dataout_18,ri_dataout_19,ri_dataout_20,ri_dataout_21,ri_dataout_22,ri_dataout_23,ri_dataout_24,ri_dataout_25,ri_dataout_26,ri_dataout_27,ri_dataout_28,ri_dataout_29,ri_dataout_30,ri_dataout_31,ri_dataout_32: std_logic;--_vector (1 to 1);
signal lo_dataout_1,lo_dataout_2,lo_dataout_3,lo_dataout_4,lo_dataout_5,lo_dataout_6,lo_dataout_7,lo_dataout_8,lo_dataout_9,lo_dataout_10,lo_dataout_11,lo_dataout_12,lo_dataout_13,lo_dataout_14,lo_dataout_15,lo_dataout_16,lo_dataout_17,lo_dataout_18,lo_dataout_19,lo_dataout_20,lo_dataout_21,lo_dataout_22,lo_dataout_23,lo_dataout_24,lo_dataout_25,lo_dataout_26,lo_dataout_27,lo_dataout_28,lo_dataout_29,lo_dataout_30,lo_dataout_31,lo_dataout_32: std_logic;--_vector (1 to 1);
signal ro_dataout_1,ro_dataout_2,ro_dataout_3,ro_dataout_4,ro_dataout_5,ro_dataout_6,ro_dataout_7,ro_dataout_8,ro_dataout_9,ro_dataout_10,ro_dataout_11,ro_dataout_12,ro_dataout_13,ro_dataout_14,ro_dataout_15,ro_dataout_16,ro_dataout_17,ro_dataout_18,ro_dataout_19,ro_dataout_20,ro_dataout_21,ro_dataout_22,ro_dataout_23,ro_dataout_24,ro_dataout_25,ro_dataout_26,ro_dataout_27,ro_dataout_28,ro_dataout_29,ro_dataout_30,ro_dataout_31,ro_dataout_32: std_logic;--_vector (1 to 1);

signal li_scanout,ri_scanout,lo_scanout,ro_scanout:  std_logic_vector(1 to 32);

component scan_ff
port (
scan_clk : in std_logic;
reset : in std_logic;
test_enable : in std_logic;
ShiftDR : in std_logic;
UpdateDR : in std_logic;
CaptureDR : in std_logic;
scan_in : in std_logic;
data_in : in std_logic;
scan_out : out std_logic;
data_out : out std_logic
);
end component;
begin

li_1<=li_in(1);
li_2<=li_in(2);
li_3<=li_in(3);
li_4<=li_in(4);
li_5<=li_in(5);
li_6<=li_in(6);
li_7<=li_in(7);
li_8<=li_in(8);
li_9<=li_in(9);
li_10<=li_in(10);
li_11<=li_in(11);
li_12<=li_in(12);
li_13<=li_in(13);
li_14<=li_in(14);
li_15<=li_in(15);
li_16<=li_in(16);
li_17<=li_in(17);
li_18<=li_in(18);
li_19<=li_in(19);
li_20<=li_in(20);
li_21<=li_in(21);
li_22<=li_in(22);
li_23<=li_in(23);
li_24<=li_in(24);
li_25<=li_in(25);
li_26<=li_in(26);
li_27<=li_in(27);
li_28<=li_in(28);
li_29<=li_in(29);
li_30<=li_in(30);
li_31<=li_in(31);
li_32<=li_in(32);

ri_1<=ri_in(1);
ri_2<=ri_in(2);
ri_3<=ri_in(3);
ri_4<=ri_in(4);
ri_5<=ri_in(5);
ri_6<=ri_in(6);
ri_7<=ri_in(7);
ri_8<=ri_in(8);
ri_9<=ri_in(9);
ri_10<=ri_in(10 );
ri_11<=ri_in(11 );
ri_12<=ri_in(12 );
ri_13<=ri_in(13 );
ri_14<=ri_in(14 );
ri_15<=ri_in(15 );
ri_16<=ri_in(16 );
ri_17<=ri_in(17 );
ri_18<=ri_in(18 );
ri_19<=ri_in(19 );
ri_20<=ri_in(20 );
ri_21<=ri_in(21 );
ri_22<=ri_in(22 );
ri_23<=ri_in(23 );
ri_24<=ri_in(24 );
ri_25<=ri_in(25 );
ri_26<=ri_in(26 );
ri_27<=ri_in(27 );
ri_28<=ri_in(28 );
ri_29<=ri_in(29 );
ri_30<=ri_in(30 );
ri_31<=ri_in(31 );
ri_32<=ri_in(32 );
lo_1<=lo_in(1);
lo_2<=lo_in(2);
lo_3<=lo_in(3);
lo_4<=lo_in(4);
lo_5<=lo_in(5);
lo_6<=lo_in(6);
lo_7<=lo_in(7);
lo_8<=lo_in(8);
lo_9<=lo_in(9);
lo_10<=lo_in(10);
lo_11<=lo_in(11);
lo_12<=lo_in(12);
lo_13<=lo_in(13);
lo_14<=lo_in(14);
lo_15<=lo_in(15);
lo_16<=lo_in(16);
lo_17<=lo_in(17);
lo_18<=lo_in(18);
lo_19<=lo_in(19);
lo_20<=lo_in(20);
lo_21<=lo_in(21);
lo_22<=lo_in(22);
lo_23<=lo_in(23);
lo_24<=lo_in(24);
lo_25<=lo_in(25);
lo_26<=lo_in(26);
lo_27<=lo_in(27);
lo_28<=lo_in(28);
lo_29<=lo_in(29);
lo_30<=lo_in(30);
lo_31<=lo_in(31);
lo_32<=lo_in(32);
ro_1<=ro_in(1);
ro_2<=ro_in(2);
ro_3<=ro_in(3);
ro_4<=ro_in(4);
ro_5<=ro_in(5);
ro_6<=ro_in(6);
ro_7<=ro_in(7);
ro_8<=ro_in(8);
ro_9<=ro_in(9);
ro_10<=ro_in(10);
ro_11<=ro_in(11);
ro_12<=ro_in(12);
ro_13<=ro_in(13);
ro_14<=ro_in(14);
ro_15<=ro_in(15);
ro_16<=ro_in(16);
ro_17<=ro_in(17);
ro_18<=ro_in(18);
ro_19<=ro_in(19);
ro_20<=ro_in(20);
ro_21<=ro_in(21);
ro_22<=ro_in(22);
ro_23<=ro_in(23);
ro_24<=ro_in(24);
ro_25<=ro_in(25);
ro_26<=ro_in(26);
ro_27<=ro_in(27);
ro_28<=ro_in(28);
ro_29<=ro_in(29);
ro_30<=ro_in(30);
ro_31<=ro_in(31);
ro_32<=ro_in(32);
ri_dataout <= ri_dataout_1 & ri_dataout_2 & ri_dataout_3 & ri_dataout_4 & ri_dataout_5 & ri_dataout_6 & ri_dataout_7 & ri_dataout_8 & ri_dataout_9 & ri_dataout_10 & ri_dataout_11 & ri_dataout_12 & ri_dataout_13 & ri_dataout_14 & ri_dataout_15 & ri_dataout_16 & ri_dataout_17 & ri_dataout_18 & ri_dataout_19 & ri_dataout_20 & ri_dataout_21 & ri_dataout_22 & ri_dataout_23 & ri_dataout_24 & ri_dataout_25 & ri_dataout_26 & ri_dataout_27 & ri_dataout_28 & ri_dataout_29 & ri_dataout_30 & ri_dataout_31 & ri_dataout_32;
ro_dataout <= ro_dataout_1 & ro_dataout_2 & ro_dataout_3 & ro_dataout_4 & ro_dataout_5 & ro_dataout_6 & ro_dataout_7 & ro_dataout_8 & ro_dataout_9 & ro_dataout_10 & ro_dataout_11 & ro_dataout_12 & ro_dataout_13 & ro_dataout_14 & ro_dataout_15 & ro_dataout_16 & ro_dataout_17 & ro_dataout_18 & ro_dataout_19 & ro_dataout_20 & ro_dataout_21 & ro_dataout_22 & ro_dataout_23 & ro_dataout_24 & ro_dataout_25 & ro_dataout_26 & ro_dataout_27 & ro_dataout_28 & ro_dataout_29 & ro_dataout_30 & ro_dataout_31 & ro_dataout_32;
lo_dataout <= lo_dataout_1 & lo_dataout_2 & lo_dataout_3 & lo_dataout_4 & lo_dataout_5 & lo_dataout_6 & lo_dataout_7 & lo_dataout_8 & lo_dataout_9 & lo_dataout_10 & lo_dataout_11 & lo_dataout_12 & lo_dataout_13 & lo_dataout_14 & lo_dataout_15 & lo_dataout_16 & lo_dataout_17 & lo_dataout_18 & lo_dataout_19 & lo_dataout_20 & lo_dataout_21 & lo_dataout_22 & lo_dataout_23 & lo_dataout_24 & lo_dataout_25 & lo_dataout_26 & lo_dataout_27 & lo_dataout_28 & lo_dataout_29 & lo_dataout_30 & lo_dataout_31 & lo_dataout_32;
li_dataout <= li_dataout_1 & li_dataout_2 & li_dataout_3 & li_dataout_4 & li_dataout_5 & li_dataout_6 & li_dataout_7 & li_dataout_8 & li_dataout_9 & li_dataout_10 & li_dataout_11 & li_dataout_12 & li_dataout_13 & li_dataout_14 & li_dataout_15 & li_dataout_16 & li_dataout_17 & li_dataout_18 & li_dataout_19 & li_dataout_20 & li_dataout_21 & li_dataout_22 & li_dataout_23 & li_dataout_24 & li_dataout_25 & li_dataout_26 & li_dataout_27 & li_dataout_28 & li_dataout_29 & li_dataout_30 & li_dataout_31 & li_dataout_32;
scan_out <= lo_scanout_32;
ri_scanout <= ri_scanout_1 & ri_scanout_2 & ri_scanout_3 & ri_scanout_4 & ri_scanout_5 & ri_scanout_6 & ri_scanout_7 & ri_scanout_8 & ri_scanout_9 & ri_scanout_10 & ri_scanout_11 & ri_scanout_12 & ri_scanout_13 & ri_scanout_14 & ri_scanout_15 & ri_scanout_16 & ri_scanout_17 & ri_scanout_18 & ri_scanout_19 & ri_scanout_20 & ri_scanout_21 & ri_scanout_22 & ri_scanout_23 & ri_scanout_24 & ri_scanout_25 & ri_scanout_26 & ri_scanout_27 & ri_scanout_28 & ri_scanout_29 & ri_scanout_30 & ri_scanout_31 & ri_scanout_32;
ro_scanout <= ro_scanout_1 & ro_scanout_2 & ro_scanout_3 & ro_scanout_4 & ro_scanout_5 & ro_scanout_6 & ro_scanout_7 & ro_scanout_8 & ro_scanout_9 & ro_scanout_10 & ro_scanout_11 & ro_scanout_12 & ro_scanout_13 & ro_scanout_14 & ro_scanout_15 & ro_scanout_16 & ro_scanout_17 & ro_scanout_18 & ro_scanout_19 & ro_scanout_20 & ro_scanout_21 & ro_scanout_22 & ro_scanout_23 & ro_scanout_24 & ro_scanout_25 & ro_scanout_26 & ro_scanout_27 & ro_scanout_28 & ro_scanout_29 & ro_scanout_30 & ro_scanout_31 & ro_scanout_32;
lo_scanout <= lo_scanout_1 & lo_scanout_2 & lo_scanout_3 & lo_scanout_4 & lo_scanout_5 & lo_scanout_6 & lo_scanout_7 & lo_scanout_8 & lo_scanout_9 & lo_scanout_10 & lo_scanout_11 & lo_scanout_12 & lo_scanout_13 & lo_scanout_14 & lo_scanout_15 & lo_scanout_16 & lo_scanout_17 & lo_scanout_18 & lo_scanout_19 & lo_scanout_20 & lo_scanout_21 & lo_scanout_22 & lo_scanout_23 & lo_scanout_24 & lo_scanout_25 & lo_scanout_26 & lo_scanout_27 & lo_scanout_28 & lo_scanout_29 & lo_scanout_30 & lo_scanout_31 & lo_scanout_32;
li_scanout <= li_scanout_1 & li_scanout_2 & li_scanout_3 & li_scanout_4 & li_scanout_5 & li_scanout_6 & li_scanout_7 & li_scanout_8 & li_scanout_9 & li_scanout_10 & li_scanout_11 & li_scanout_12 & li_scanout_13 & li_scanout_14 & li_scanout_15 & li_scanout_16 & li_scanout_17 & li_scanout_18 & li_scanout_19 & li_scanout_20 & li_scanout_21 & li_scanout_22 & li_scanout_23 & li_scanout_24 & li_scanout_25 & li_scanout_26 & li_scanout_27 & li_scanout_28 & li_scanout_29 & li_scanout_30 & li_scanout_31 & li_scanout_32;
scan_ff1: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => scan_in, data_in =>li_1, scan_out => li_scanout_1,data_out => li_dataout_1); 
scan_ff2: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_1, data_in =>li_2, scan_out => li_scanout_2,data_out => li_dataout_2);
scan_ff3: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_2, data_in =>li_3, scan_out => li_scanout_3,data_out => li_dataout_3);
scan_ff4: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_3, data_in =>li_4, scan_out => li_scanout_4,data_out => li_dataout_4);
scan_ff5: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_4, data_in =>li_5, scan_out => li_scanout_5,data_out => li_dataout_5);
scan_ff6: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_5, data_in =>li_6, scan_out => li_scanout_6,data_out => li_dataout_6);
scan_ff7: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_6, data_in =>li_7, scan_out => li_scanout_7,data_out => li_dataout_7);
scan_ff8: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_7, data_in =>li_8, scan_out => li_scanout_8,data_out => li_dataout_8);
scan_ff9: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_8, data_in =>li_9, scan_out => li_scanout_9,data_out => li_dataout_9);
scan_ff10: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_9, data_in =>li_10, scan_out => li_scanout_10,data_out => li_dataout_10);
scan_ff11: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_10, data_in =>li_11, scan_out => li_scanout_11,data_out => li_dataout_11);
scan_ff12: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_11, data_in =>li_12, scan_out => li_scanout_12,data_out => li_dataout_12);
scan_ff13: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_12, data_in =>li_13, scan_out => li_scanout_13,data_out => li_dataout_13);
scan_ff14: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_13, data_in =>li_14, scan_out => li_scanout_14,data_out => li_dataout_14);
scan_ff15: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_14, data_in =>li_15, scan_out => li_scanout_15,data_out => li_dataout_15);
scan_ff16: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_15, data_in =>li_16, scan_out => li_scanout_16,data_out => li_dataout_16);
scan_ff17: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_16, data_in =>li_17, scan_out => li_scanout_17,data_out => li_dataout_17);
scan_ff18: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_17, data_in =>li_18, scan_out => li_scanout_18,data_out => li_dataout_18);
scan_ff19: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_18, data_in =>li_19, scan_out => li_scanout_19,data_out => li_dataout_19);
scan_ff20: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_19, data_in =>li_20, scan_out => li_scanout_20,data_out => li_dataout_20);
scan_ff21: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_20, data_in =>li_21, scan_out => li_scanout_21,data_out => li_dataout_21);
scan_ff22: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_21, data_in =>li_22, scan_out => li_scanout_22,data_out => li_dataout_22);
scan_ff23: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_22, data_in =>li_23, scan_out => li_scanout_23,data_out => li_dataout_23);
scan_ff24: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_23, data_in =>li_24, scan_out => li_scanout_24,data_out => li_dataout_24);
scan_ff25: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_24, data_in =>li_25, scan_out => li_scanout_25,data_out => li_dataout_25);
scan_ff26: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_25, data_in =>li_26, scan_out => li_scanout_26,data_out => li_dataout_26);
scan_ff27: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_26, data_in =>li_27, scan_out => li_scanout_27,data_out => li_dataout_27);
scan_ff28: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_27, data_in =>li_28, scan_out => li_scanout_28,data_out => li_dataout_28);
scan_ff29: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_28, data_in =>li_29, scan_out => li_scanout_29,data_out => li_dataout_29);
scan_ff30: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_29, data_in =>li_30, scan_out => li_scanout_30,data_out => li_dataout_30);
scan_ff31: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_30, data_in =>li_31, scan_out => li_scanout_31,data_out => li_dataout_31);
scan_ff32: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_31, data_in =>li_32, scan_out => li_scanout_32,data_out => li_dataout_32);

scan_ff33: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => li_scanout_32, data_in =>ri_1, scan_out => ri_scanout_1,data_out => ri_dataout_1);
scan_ff34: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_1, data_in =>ri_2, scan_out => ri_scanout_2,data_out => ri_dataout_2);
scan_ff35: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_2, data_in =>ri_3, scan_out => ri_scanout_3,data_out => ri_dataout_3);
scan_ff36: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_3, data_in =>ri_4, scan_out => ri_scanout_4,data_out => ri_dataout_4);
scan_ff37: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_4, data_in =>ri_5, scan_out => ri_scanout_5,data_out => ri_dataout_5);
scan_ff38: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_5, data_in =>ri_6, scan_out => ri_scanout_6,data_out => ri_dataout_6);
scan_ff39: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_6, data_in =>ri_7, scan_out => ri_scanout_7,data_out => ri_dataout_7);
scan_ff40: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_7, data_in =>ri_8, scan_out => ri_scanout_8,data_out => ri_dataout_8);
scan_ff41: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_8, data_in =>ri_9, scan_out => ri_scanout_9,data_out => ri_dataout_9);
scan_ff42: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_9, data_in =>ri_10, scan_out => ri_scanout_10,data_out => ri_dataout_10);
scan_ff43: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_10, data_in =>ri_11, scan_out => ri_scanout_11,data_out => ri_dataout_11);
scan_ff44: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_11, data_in =>ri_12, scan_out => ri_scanout_12,data_out => ri_dataout_12);
scan_ff45: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_12, data_in =>ri_13, scan_out => ri_scanout_13,data_out => ri_dataout_13);
scan_ff46: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_13, data_in =>ri_14, scan_out => ri_scanout_14,data_out => ri_dataout_14);
scan_ff47: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_14, data_in =>ri_15, scan_out => ri_scanout_15,data_out => ri_dataout_15);
scan_ff48: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_15, data_in =>ri_16, scan_out => ri_scanout_16,data_out => ri_dataout_16);
scan_ff49: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_16, data_in =>ri_17, scan_out => ri_scanout_17,data_out => ri_dataout_17);
scan_ff50: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_17, data_in =>ri_18, scan_out => ri_scanout_18,data_out => ri_dataout_18);
scan_ff51: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_18, data_in =>ri_19, scan_out => ri_scanout_19,data_out => ri_dataout_19);
scan_ff52: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_19, data_in =>ri_20, scan_out => ri_scanout_20,data_out => ri_dataout_20);
scan_ff53: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_20, data_in =>ri_21, scan_out => ri_scanout_21,data_out => ri_dataout_21);
scan_ff54: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_21, data_in =>ri_22, scan_out => ri_scanout_22,data_out => ri_dataout_22);
scan_ff55: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_22, data_in =>ri_23, scan_out => ri_scanout_23,data_out => ri_dataout_23);
scan_ff56: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_23, data_in =>ri_24, scan_out => ri_scanout_24,data_out => ri_dataout_24);
scan_ff57: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_24, data_in =>ri_25, scan_out => ri_scanout_25,data_out => ri_dataout_25);
scan_ff58: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_25, data_in =>ri_26, scan_out => ri_scanout_26,data_out => ri_dataout_26);
scan_ff59: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_26, data_in =>ri_27, scan_out => ri_scanout_27,data_out => ri_dataout_27);
scan_ff60: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_27, data_in =>ri_28, scan_out => ri_scanout_28,data_out => ri_dataout_28);
scan_ff61: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_28, data_in =>ri_29, scan_out => ri_scanout_29,data_out => ri_dataout_29);
scan_ff62: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_29, data_in =>ri_30, scan_out => ri_scanout_30,data_out => ri_dataout_30);
scan_ff63: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_30, data_in =>ri_31, scan_out => ri_scanout_31,data_out => ri_dataout_31);
scan_ff64: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_31, data_in =>ri_32, scan_out => ri_scanout_32,data_out => ri_dataout_32);

scan_ff65: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ri_scanout_32, data_in =>ro_1, scan_out => ro_scanout_1,data_out => ro_dataout_1);
scan_ff66: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_1, data_in =>ro_2, scan_out => ro_scanout_2,data_out => ro_dataout_2);
scan_ff67: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_2, data_in =>ro_3, scan_out => ro_scanout_3,data_out => ro_dataout_3);
scan_ff68: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_3, data_in =>ro_4, scan_out => ro_scanout_4,data_out => ro_dataout_4);
scan_ff69: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_4, data_in =>ro_5, scan_out => ro_scanout_5,data_out => ro_dataout_5);
scan_ff70: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_5, data_in =>ro_6, scan_out => ro_scanout_6,data_out => ro_dataout_6);
scan_ff71: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_6, data_in =>ro_7, scan_out => ro_scanout_7,data_out => ro_dataout_7);
scan_ff72: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_7, data_in =>ro_8, scan_out => ro_scanout_8,data_out => ro_dataout_8);
scan_ff73: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_8, data_in =>ro_9, scan_out => ro_scanout_9,data_out => ro_dataout_9);
scan_ff74: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_9, data_in =>ro_10, scan_out => ro_scanout_10,data_out => ro_dataout_10);
scan_ff75: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_10, data_in =>ro_11, scan_out => ro_scanout_11,data_out => ro_dataout_11);
scan_ff76: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_11, data_in =>ro_12, scan_out => ro_scanout_12,data_out => ro_dataout_12);
scan_ff77: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_12, data_in =>ro_13, scan_out => ro_scanout_13,data_out => ro_dataout_13);
scan_ff78: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_13, data_in =>ro_14, scan_out => ro_scanout_14,data_out => ro_dataout_14);
scan_ff79: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_14, data_in =>ro_15, scan_out => ro_scanout_15,data_out => ro_dataout_15);
scan_ff80: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_15, data_in =>ro_16, scan_out => ro_scanout_16,data_out => ro_dataout_16);
scan_ff81: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_16, data_in =>ro_17, scan_out => ro_scanout_17,data_out => ro_dataout_17);
scan_ff82: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_17, data_in =>ro_18, scan_out => ro_scanout_18,data_out => ro_dataout_18);
scan_ff83: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_18, data_in =>ro_19, scan_out => ro_scanout_19,data_out => ro_dataout_19);
scan_ff84: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_19, data_in =>ro_20, scan_out => ro_scanout_20,data_out => ro_dataout_20);
scan_ff85: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_20, data_in =>ro_21, scan_out => ro_scanout_21,data_out => ro_dataout_21);
scan_ff86: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_21, data_in =>ro_22, scan_out => ro_scanout_22,data_out => ro_dataout_22);
scan_ff87: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_22, data_in =>ro_23, scan_out => ro_scanout_23,data_out => ro_dataout_23);
scan_ff88: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_23, data_in =>ro_24, scan_out => ro_scanout_24,data_out => ro_dataout_24);
scan_ff89: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_24, data_in =>ro_25, scan_out => ro_scanout_25,data_out => ro_dataout_25);
scan_ff90: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_25, data_in =>ro_26, scan_out => ro_scanout_26,data_out => ro_dataout_26);
scan_ff91: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_26, data_in =>ro_27, scan_out => ro_scanout_27,data_out => ro_dataout_27);
scan_ff92: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_27, data_in =>ro_28, scan_out => ro_scanout_28,data_out => ro_dataout_28);
scan_ff93: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_28, data_in =>ro_29, scan_out => ro_scanout_29,data_out => ro_dataout_29);
scan_ff94: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_29, data_in =>ro_30, scan_out => ro_scanout_30,data_out => ro_dataout_30);
scan_ff95: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_30, data_in =>ro_31, scan_out => ro_scanout_31,data_out => ro_dataout_31);
scan_ff96: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_31, data_in =>ro_32, scan_out => ro_scanout_32,data_out => ro_dataout_32);

scan_ff97: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => ro_scanout_32, data_in =>lo_1, scan_out => lo_scanout_1,data_out => lo_dataout_1);
scan_ff98: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_1, data_in =>lo_2, scan_out => lo_scanout_2,data_out => lo_dataout_2);
scan_ff99: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_2, data_in =>lo_3, scan_out => lo_scanout_3,data_out => lo_dataout_3);
scan_ff100: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_3, data_in =>lo_4, scan_out => lo_scanout_4,data_out => lo_dataout_4);
scan_ff101: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_4, data_in =>lo_5, scan_out => lo_scanout_5,data_out => lo_dataout_5);
scan_ff102: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_5, data_in =>lo_6, scan_out => lo_scanout_6,data_out => lo_dataout_6);
scan_ff103: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_6, data_in =>lo_7, scan_out => lo_scanout_7,data_out => lo_dataout_7);
scan_ff104: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_7, data_in =>lo_8, scan_out => lo_scanout_8,data_out => lo_dataout_8);
scan_ff105: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_8, data_in =>lo_9, scan_out => lo_scanout_9,data_out => lo_dataout_9);
scan_ff106: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_9, data_in =>lo_10, scan_out => lo_scanout_10,data_out => lo_dataout_10);
scan_ff107: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_10, data_in =>lo_11, scan_out => lo_scanout_11,data_out => lo_dataout_11);
scan_ff108: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_11, data_in =>lo_12, scan_out => lo_scanout_12,data_out => lo_dataout_12);
scan_ff109: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_12, data_in =>lo_13, scan_out => lo_scanout_13,data_out => lo_dataout_13);
scan_ff110: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_13, data_in =>lo_14, scan_out => lo_scanout_14,data_out => lo_dataout_14);
scan_ff111: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_14, data_in =>lo_15, scan_out => lo_scanout_15,data_out => lo_dataout_15);
scan_ff112: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_15, data_in =>lo_16, scan_out => lo_scanout_16,data_out => lo_dataout_16);
scan_ff113: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_16, data_in =>lo_17, scan_out => lo_scanout_17,data_out => lo_dataout_17);
scan_ff114: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_17, data_in =>lo_18, scan_out => lo_scanout_18,data_out => lo_dataout_18);
scan_ff115: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_18, data_in =>lo_19, scan_out => lo_scanout_19,data_out => lo_dataout_19);
scan_ff116: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_19, data_in =>lo_20, scan_out => lo_scanout_20,data_out => lo_dataout_20);
scan_ff117: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_20, data_in =>lo_21, scan_out => lo_scanout_21,data_out => lo_dataout_21);
scan_ff118: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_21, data_in =>lo_22, scan_out => lo_scanout_22,data_out => lo_dataout_22);
scan_ff119: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_22, data_in =>lo_23, scan_out => lo_scanout_23,data_out => lo_dataout_23);
scan_ff120: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_23, data_in =>lo_24, scan_out => lo_scanout_24,data_out => lo_dataout_24);
scan_ff121: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_24, data_in =>lo_25, scan_out => lo_scanout_25,data_out => lo_dataout_25);
scan_ff122: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_25, data_in =>lo_26, scan_out => lo_scanout_26,data_out => lo_dataout_26);
scan_ff123: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_26, data_in =>lo_27, scan_out => lo_scanout_27,data_out => lo_dataout_27);
scan_ff124: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_27, data_in =>lo_28, scan_out => lo_scanout_28,data_out => lo_dataout_28);
scan_ff125: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_28, data_in =>lo_29, scan_out => lo_scanout_29,data_out => lo_dataout_29);
scan_ff126: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_29, data_in =>lo_30, scan_out => lo_scanout_30,data_out => lo_dataout_30);
scan_ff127: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_30, data_in =>lo_31, scan_out => lo_scanout_31,data_out => lo_dataout_31);
scan_ff128: scan_ff port map(scan_clk => scan_clk,CaptureDR=>CaptureDR,UpdateDR=>UpdateDR,ShiftDR=>ShiftDR,  reset => reset, test_enable => test_enable, scan_in => lo_scanout_31, data_in =>lo_32, scan_out => lo_scanout_32,data_out => lo_dataout_32);



end behaviour;