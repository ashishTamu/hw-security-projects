module FeistelNetwork()

endmodule
