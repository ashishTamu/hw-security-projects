module InitialPermutation();
endmodule
