module RoundOperation()
endmodule
