module FinalPermutation()
endmodule
