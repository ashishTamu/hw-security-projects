module Decryption()
endmodule
