module RoundKeyGenerator()

endmodule

