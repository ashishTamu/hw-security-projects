/* 
 * Feistal Function SBOX Permutation
 * for DES encryption algorithm
 * 
 */

module SBox(wOutputData, wInputData);
   
   //input is 48 bit
   input wire [47:0] wInputData ;
   //output is 32 bit
   output wire [31:0] wOutputData ;


   
endmodule // SBox

