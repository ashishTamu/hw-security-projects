module InitialPermutation();
   
endmodule // InitialPermutation

