module KeyExpansionPermChoice2(wOutputData, wInputData);


   input wire [47:0] wInputData ;

   output wire [47:0] wOutputData ;
endmodule // KeyExpansionPermChoice2
