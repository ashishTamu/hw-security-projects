module KeyExpansionPermChoice1(wOutputData, wInputData);

   //input is 32 bit
   input wire [31:0] wInputData ;
   //output is 32 bit
   output wire [31:0] wOutputData ;
endmodule // KeyExpansionPermChoice1
