module ExpansionBox()
endmodule
