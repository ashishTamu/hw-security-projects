module InitialPermutation();
endmodule // InitialPermutation
