module SBox()
endmodule
