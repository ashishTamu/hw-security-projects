module Decryption();
   
endmodule // Decryption

